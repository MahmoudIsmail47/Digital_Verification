module RAM_tb_A1 ();





endmodule